module test ( input T,R, // Мы создаем Счетчик, по аналогии с теорией, создаем D триггер и к нему комбинационную схему. Нам необходимо получить T триггер и комбинационку к нему
              input C,
              output [23:0]Q);
        
         wire [23:0] Y = {24{!R}} & ({24{T}} & (Q + 1'd1) |  ({24{!T}} & Q)); /* Это описание комбинационной схемы для того, чтобы получить счетчик в итоге. Если T=1, то выражение T & (Q + 1d'1)
                                                        позволяет производить счет, получается Q+1. А выражение (!T & Q) дает по сути 0.
                                                        Если T=1, то выражение T & (Q + 1d'1) уже не работает и выдает 0, а (!T & Q) дает нам хранение предыдущего состояния 
                                                        R - сброс, мы сделаем хитрый способ вставить сюда сброс. Сделаем R инверсным, получится, если сброс в 1, то все наши 
                                                        выражения в скобках не работают. Если R будет = 0, то выражение работает  
                                                        Еще мы не можем оставлять R и T в одноразрядном значении (т.к у нас 24 разряда), поэтому прибегнем к конкатенации{} 
                                                        Компилятор каким-то образом пониает что такое 1'd1.*/
                                        
         DT DT [23:0] (.q(Q), .D(Y), .C(C));    // Это у нас массив модулей D триггера (этот модуль описан ниже)
endmodule

module DT(input D, input C, output Q);
	    DFF DT (
				.d(D),         // Это по сути наши данные в D триггер 
				.clk(C),       // Это clk, наш тактовый сигнал для D Триггера
				.clrn(1'd1),   // Это Асинхронный сброс, он нам не нужен, поэтому ставим 1, так как инверсия
				.prn(1'd1),    // Это асинхронный вход установки (тоже нам не нужен и тоже инверсный)
				.q(Q)          // Ну а это логично - выход
				);
endmodule



/* Этот код по сути показывает нам внутреннее состояние. Но нам необходимо это перенести на плату, поэтому я сделаю вторую часть кода, в котором произойдут некоторые изменения