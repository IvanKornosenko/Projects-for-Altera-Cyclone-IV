library verilog;
use verilog.vl_types.all;
entity sev_seg_tb is
end sev_seg_tb;
