module test ( (* chip_pin = "88" *)input nT, // Вторая часть, пытаемся реализовать на плате. nT и nR означают, что мы должны подавать их инверсными, потому что кнопка на плате дает "0" при нажатии
              (* chip_pin = "89" *)input nR,
              (* chip_pin = "23" *)input C,
              (* chip_pin = "87" *)output LedQ); //Делаем обозначение вывода на светодиод. Выводить будем 23-й разряд, т.е. старший. 
        wire [23:0] Q;
        wire TQ, RQ; // nT и nR проинвертировали и они стали TQ и RQ
        DT Sync [1:0] (.Q({TQ, RQ}), .D({!nT, !nR}), .C(C)); /* Нам нужно засинхронизировать R и T, потому что мы будем подавать их с кнопки. Кнопку мы будем нажимать 
                                                                асинхронно тактовому сигналу. Для этой синхронизации используем шаблон D триггера */
        wire [23:0] Y = {24{!RQ}} & ({24{TQ}} & (Q + 1'd1) |  ({24{!TQ}} & Q)); // T заменяем на TQ, а R заменяем на RQ.
                                        
        DT DT [23:0] (.Q(Q), .D(Y), .C(C));    
        assign LedQ = !Q[23]; // Наблюдаем за 23 разрядом (Диод кстати тоже инвертировали, потому что он по умолчанию в 1)
endmodule

module DT(input D, input C, output Q);
	    DFF DT (
				.d(D),         // Это по сути наши данные в D триггер 
				.clk(C),       // Это clk, наш тактовый сигнал для D Триггера
				.clrn(1'd1),   // Это Асинхронный сброс, он нам не нужен, поэтому ставим 1, так как инверсия
				.prn(1'd1),    // Это асинхронный вход установки (тоже нам не нужен и тоже инверсный)
				.q(Q)          // Ну а это логично - выход
				);
endmodule

