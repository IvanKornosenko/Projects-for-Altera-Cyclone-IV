module sev_seg_top (
    input CLOCK_50,             //50 МГц, это тактовый сигнал на самой плате
    input [1:0] KEY,            //нажатие кнопки
    output [6:0] HEX0,          //вывод на сегменты g f e d c b a (На моей плате семигегментник один, с общими выводами на 4 разряда )
    output DIG4                 //вывод на 4-й разряд

);
    reg [26:0] cnt;             /*это счетчтик, делитель частоты. Мы будем делить тактовый сигнал. Внутри модуля мы создаем 2 регистра
                                 cnt - 27 бит (может считать до 134 миллионов), он нужен, чтобы из 50 МГц сделать 1 Гц
                                 digit - 4 бита, чтобы отображать числа от 0 до 15 на семисегментниках*/
    reg [3:0] digit;
    always @(posedge CLOCK_50 or negedge KEY[0])
    begin
        if (!KEY[0])            //Если кнопка нажата (KEY[0] = 0)
        begin
        cnt <=0;                //обнуляем счетчик
        digit <=0;              //и цифру тоже
        end
            else                //иначе, если кнопка не нажата
            begin   
                if (cnt == 27'd49_999_999) //если счетчик достигнет 49 999 999
                begin
                    cnt <= 0;               //обнуляем счетчик
                    digit <= digit + 1;     //и увеличиваем цифру
                end
                    else                    //иначе
                        begin
                        cnt <= cnt + 1;     //просто считаем дальше
                        end
            end
    end     
   /*По сути получается, что 50 МГц = 50 000 000 тактов в секунду
   Мы считаем до 49999999, это почти ровно 1 секунда.
   Когда дошли, обгуляем счетчик и увеличиваем цифру
   Цифра меняется раз в секунду */

   //Подключаем декодер
   sev_seg u_hex0 (
    .digit(digit),
    .segments(HEX0)
   );

   //включаем только один 4-й разряд на плате
   assign DIG4 = 1'b0;              //0 - это у нас "включено"
endmodule
